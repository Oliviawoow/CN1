// CN1 -  schelet lab02

module modul02(
  output out,
  input in
  );

  assign out = ~in;

endmodule
